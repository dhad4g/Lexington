`timescale 1ns/1ps

`include "axi4_lite.sv"


module axi4_lite_crossbar_TB;

    

endmodule
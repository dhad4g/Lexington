`timescale 1ns/1ps

`include "rv32.sv"
`include "saratoga.sv"
import saratoga::*;


module decoder (
        // clock not needed; module is purely combinatorial
        // reset not needed; module is stateless

        input  rv32::word inst,                     // instruction bits from fetch
        input  rv32::word pc,                       // current program counter
        output logic branch,                        // jump/branch taken
        output rv32::word branch_addr,              // next PC calculation

        // Register File Ports
        output logic rs1_en,                        // register source 1 enable
        output rv32::gpr_addr_t rs1_addr,           // register source 1 address
        input  rv32::word rs1_data,                 // register source 1 data
        output logic rs2_en,                        // register source 2 enable
        output rv32::gpr_addr_t rs2_addr,           // register source 2 address
        input  rv32::word rs2_data,                 // register source 2 data

        // CSR Ports
        output logic csr_rd_en,                     // CSR read enable
        output logic csr_explicit_rd,               // CSR explicit read flag
        output rv32::csr_addr_t csr_addr,           // CSR read address
        input  rv32::word csr_rd_data,              // CSR read data
        input logic csr_addr_is_atomic,             // indicates CSR is atomic
        input logic csr_addr_is_illegal,            // indicates CSR does not exists or incorrect permission
        output logic atomic_csr,                    // indicates atomic CSR write

        // ALU Ports
        output alu_op_t alu_op,                     // ALU operation select
        output rv32::word src1,                     // ALU left-side operand
        output rv32::word src2,                     // ALU right-side operand

        // Load/Store Ports
        output lsu_op_t lsu_op,                     // LSU operation select
        output rv32::word alt_data,                 // LSU alternate data
        output rv32::gpr_addr_t dest_addr,          // LSU destination register address

        // Exception Flags
        output logic illegal_inst,                  // illegal instruction flag
        output logic inst_misaligned,               // instruction misaligned flag, generated by jump/branch instruction
        output logic ecall,                         // environment call exception flag
        output logic ebreak,                        // environment breakpoint exception flag
        output logic mret                           // MRET instruction flag
    );

    localparam OPCODE_WIDTH  = 7;   // RISC-V major opcode width

    // Major OpCode Values
    localparam OP       = 7'b011_0011;
    localparam OP_IMM   = 7'b001_0011;
    localparam LUI      = 7'b011_0111;
    localparam AUIPC    = 7'b001_0111;
    localparam JAL      = 7'b110_1111;
    localparam JALR     = 7'b110_0111;
    localparam BRANCH   = 7'b110_0011;
    localparam LOAD     = 7'b000_0011;
    localparam STORE    = 7'b010_0011;
    localparam MISC_MEM = 7'b000_1111;
    localparam SYSTEM   = 7'b111_0011;

    // Funct7 and Funct3 Field Values
    localparam FUNCT7_ZERO      = 7'b000_0000;
    localparam FUNCT7_BIT30     = 7'b010_0000;
    // arithmetic and logic instructions funct3
    localparam FUNCT3_ADD_SUB   = 3'b000;
    localparam FUNCT3_SHIFT_L   = 3'b001;
    localparam FUNCT3_SLT       = 3'b010;
    localparam FUNCT3_SLTU      = 3'b011;
    localparam FUNCT3_XOR       = 3'b100;
    localparam FUNCT3_SHIFT_R   = 3'b101;
    localparam FUNCT3_OR        = 3'b110;
    localparam FUNCT3_AND       = 3'b111;
    // branch instructions funct3
    localparam FUNCT3_BEQ       = 3'b000;
    localparam FUNCT3_BNE       = 3'b001;
    localparam FUNCT3_BLT       = 3'b100;
    localparam FUNCT3_BGE       = 3'b101;
    localparam FUNCT3_BLTU      = 3'b110;
    localparam FUNCT3_BGEU      = 3'b111;
    // load/store instruction funct3
    localparam FUNCT3_LB        = 3'b000;
    localparam FUNCT3_LH        = 3'b001;
    localparam FUNCT3_LW        = 3'b010;
    localparam FUNCT3_LBU       = 3'b100;
    localparam FUNCT3_LHU       = 3'b101;
    localparam FUNCT3_SB        = 3'b000;
    localparam FUNCT3_SH        = 3'b001;
    localparam FUNCT3_SW        = 3'b010;
    // fence instruction funct3
    localparam FUNCT3_FENCE     = 3'b000;
    localparam FUNCT3_FENCE_I   = 3'b001;
    // CSR instruction funct3
    localparam FUNCT3_CSRRW     = 3'b001;
    localparam FUNCT3_CSRRS     = 3'b010;
    localparam FUNCT3_CSRRC     = 3'b011;
    localparam FUNCT3_CSRRWI    = 3'b101;
    localparam FUNCT3_CSRRSI    = 3'b110;
    localparam FUNCT3_CSRRCI    = 3'b111;
    // system instructions funct12
    localparam FUNCT12_ECALL    = 12'b0000_0000_0000;
    localparam FUNCT12_EBREAK   = 12'b0000_0000_0001;
    localparam FUNCT12_MRET     = 12'b0011_0000_0010;
    localparam FUNCT12_WFI      = 12'b0001_0000_0101;


    // RISC-V instruction fields
    logic [OPCODE_WIDTH-1:0] opcode;
    logic [2:0] funct3;
    logic [6:0] funct7;
    logic [11:0] funct12;
    assign opcode       = inst[6:0];
    assign dest_addr    = inst[11:7];   // output port
    assign funct3       = inst[14:12];
    assign rs1_addr     = inst[19:15];  // output port
    assign rs2_addr     = inst[24:20];  // output port
    assign funct7       = inst[31:25];
    assign funct12      = inst[31:20];
    assign csr_addr     = inst[31:20];  // output port

    assign inst_misaligned = (|branch_addr[1:0]) & branch;

    // Internal signed variants
    rv32::signed_word _src1;
    rv32::signed_word _src2;
    assign _src1 = src1;
    assign _src2 = src2;

    // Decode immediate value
    logic [31:0] immediate;
    always_comb begin
        case (opcode)
            OP_IMM:     immediate = { {20{inst[31]}}, inst[31:20] }; // sign-extended 12-bit imm[11:0]
            LUI, AUIPC: immediate = { inst[31:12], {12{1'b0}} }; // 20-bit upper-immediate imm[31:12], lower bits zero filled
            JAL:        immediate = { {12{inst[31]}}, inst[19:12], inst[20], inst[30:21], 1'b0 }; // sign-extended 20-bit imm[20:1], lowest bit zeroed
            JALR:       immediate = { {20{inst[31]}}, inst[31:20] }; // sign-extended 12-bit imm[11:0]
            BRANCH:     immediate = { {20{inst[31]}}, inst[7], inst[30:25], inst[11:8], 1'b0 }; // signed-extended 12-bit imm[12:1], lowest bit zeroed
            LOAD:       immediate = { {20{inst[31]}}, inst[31:20] }; // sign-extended 12-bit imm[11:0]
            STORE:      immediate = { {20{inst[31]}}, inst[31:25], inst[11:7] }; // sign-extended 12-bit imm[11:0]
            MISC_MEM:   immediate = { {20{inst[31]}}, inst[31:20] }; // sign-extended 12-bit imm[11:0]
            default:    immediate = { {20{inst[31]}}, inst[31:20] }; // most common decoding as default
        endcase
    end

    always_comb begin
        // defaults for exception flags, overwrite per instruction
        atomic_csr = 0;
        illegal_inst = 0;
        ecall = 0;
        ebreak = 0;
        mret = 0;
        case (opcode)

            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: OP Instructions
            ////////////////////////////////////////////////////////////
            OP: begin
                branch = 0;
                branch_addr = 0;
                // Source read enable
                rs1_en = 1;
                rs2_en = 1;
                csr_rd_en = 0;
                csr_explicit_rd = 0;
                // Source and alt data
                src1 = rs1_data;
                src2 = rs2_data;
                alt_data = 0;
                // LSU OP
                lsu_op = LSU_REG;
                // ALU OP
                if (funct7 == FUNCT7_ZERO) begin
                    case (funct3)
                        FUNCT3_ADD_SUB: alu_op = ALU_ADD;
                        FUNCT3_SHIFT_L: alu_op = ALU_SLL;
                        FUNCT3_SLT:     alu_op = ALU_SLT;
                        FUNCT3_SLTU:    alu_op = ALU_SLTU;
                        FUNCT3_XOR:     alu_op = ALU_XOR;
                        FUNCT3_SHIFT_R: alu_op = ALU_SRL;
                        FUNCT3_OR:      alu_op = ALU_OR;
                        FUNCT3_AND:     alu_op = ALU_AND;
                        default: begin
                            alu_op = ALU_NOP;
                            lsu_op = LSU_NOP;
                            illegal_inst = 1;
                        end
                    endcase
                end
                else if (funct7 == FUNCT7_BIT30) begin
                    case (funct3)
                        FUNCT3_ADD_SUB: alu_op = ALU_SUB;
                        FUNCT3_SHIFT_R: alu_op = ALU_SRA;
                        default: begin
                            alu_op = ALU_NOP;
                            lsu_op = LSU_NOP;
                            illegal_inst = 1;
                        end
                    endcase
                end
                else begin
                    alu_op = ALU_NOP;
                    lsu_op = LSU_NOP;
                    illegal_inst = 1;
                end
            end
            ////////////////////////////////////////////////////////////
            // END: OP Instructions
            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: OP-IMM Instructions
            ////////////////////////////////////////////////////////////
            OP_IMM: begin
                branch          = 0;
                branch_addr     = 0;
                rs1_en          = 1;
                rs2_en          = 0;
                csr_rd_en       = 0;
                csr_explicit_rd = 0;
                src1            = rs1_data;
                src2            = immediate;
                alt_data        = 0;
                lsu_op          = LSU_REG;
                // ALU OP
                case (funct3)
                    FUNCT3_ADD_SUB: alu_op = ALU_ADD;
                    FUNCT3_SHIFT_L: alu_op = ALU_SLL;
                    FUNCT3_SLT:     alu_op = ALU_SLT;
                    FUNCT3_SLTU:    alu_op = ALU_SLTU;
                    FUNCT3_XOR:     alu_op = ALU_XOR;
                    FUNCT3_SHIFT_R: alu_op = ALU_SRL;
                    FUNCT3_OR:      alu_op = ALU_OR;
                    FUNCT3_AND:     alu_op = ALU_AND;
                    default:
                        begin
                            alu_op = ALU_NOP;
                            lsu_op = LSU_NOP;
                            illegal_inst = 1;
                        end
                endcase
            end
            ////////////////////////////////////////////////////////////
            // END: OP-IMM Instructions
            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: LUI/AUIPC Instructions
            ////////////////////////////////////////////////////////////
            LUI, AUIPC: begin
                branch          = 0;
                branch_addr     = 0;
                rs1_en          = 0;
                rs2_en          = 0;
                csr_rd_en       = 0;
                csr_explicit_rd = 0;
                src1            = (opcode == AUIPC) ? pc : 0;
                src2            = immediate;
                alt_data        = 0;
                alu_op          = ALU_ADD;
                lsu_op          = LSU_REG;
            end
            ////////////////////////////////////////////////////////////
            // END: LUI/AUIPC Instructions
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: JAL/JALR Instruction
            ////////////////////////////////////////////////////////////
            JAL, JALR: begin
                branch          = 1;
                rs1_en          = (opcode == JALR) ? 1 : 0;
                rs2_en          = 0;
                csr_rd_en       = 0;
                csr_explicit_rd = 0;
                src1            = pc;
                src2            = 4;
                alt_data        = 0;
                alu_op          = ALU_ADD;
                lsu_op          = LSU_REG;
                // calculate jump address
                if (opcode == JAL) begin
                    branch_addr = pc + immediate;
                end
                else begin // JALR
                    // sign-extended immediate, lowest bit zeroed after calculation
                    branch_addr[31:1] = (rs1_data + immediate) >> 1;
                    branch_addr[0]    = 0;
                end
                if (inst_misaligned) begin
                    lsu_op = LSU_NOP;
                end
            end
            ////////////////////////////////////////////////////////////
            // END: JAL/JALR Instruction
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: BRANCH Instructions
            ////////////////////////////////////////////////////////////
            BRANCH: begin
                rs1_en          = 1;
                rs2_en          = 1;
                csr_rd_en       = 0;
                csr_explicit_rd = 0;
                src1            = rs1_data;
                src2            = rs2_data;
                alt_data        = 0;
                alu_op          = ALU_NOP;
                lsu_op          = LSU_NOP;
                // Branch address calculation
                // sign-extended immediate, lowest bit zero
                branch_addr     = pc + immediate;
                // Branch condition
                case (funct3)
                    FUNCT3_BEQ:     branch = (_src1 == _src2);  // branch if equal
                    FUNCT3_BNE:     branch = (_src1 != _src2);  // branch if not equal
                    FUNCT3_BLT:     branch = (_src1 <  _src2);  // branch if less than
                    FUNCT3_BGE:     branch = (_src1 >= _src2);  // branch if greater than or equal
                    FUNCT3_BLTU:    branch = (src1 <  src2);  // branch if less than unsigned
                    FUNCT3_BGEU:    branch = (src1 >= src2);  // branch if greater than or equal unsigned
                    default: begin
                        branch  = 0;
                        illegal_inst = 1;
                    end
                endcase
            end
            ////////////////////////////////////////////////////////////
            // END: BRANCH Instructions
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: LOAD/STORE Instructions
            ////////////////////////////////////////////////////////////
            LOAD, STORE: begin
                branch          = 0;
                branch_addr     = 0;
                rs1_en          = 1;
                rs2_en          = (opcode == STORE) ? 1 : 0;
                csr_rd_en       = 0;
                csr_explicit_rd = 0;
                src1            = rs1_data;
                src2            = immediate;
                alt_data        = (opcode == STORE) ? rs2_data : 0;
                alu_op          = ALU_ADD;
                if (opcode == LOAD) begin
                    case (funct3)
                        FUNCT3_LB:  lsu_op = LSU_LB;
                        FUNCT3_LH:  lsu_op = LSU_LH;
                        FUNCT3_LW:  lsu_op = LSU_LW;
                        FUNCT3_LBU: lsu_op = LSU_LBU;
                        FUNCT3_LHU: lsu_op = LSU_LHU;
                        default: begin
                            lsu_op = LSU_NOP;
                            illegal_inst = 1;
                        end
                    endcase
                end
                else begin // STORE
                    case (funct3)
                        FUNCT3_SB:  lsu_op = LSU_SB;
                        FUNCT3_SH:  lsu_op = LSU_SH;
                        FUNCT3_SW:  lsu_op = LSU_SW;
                        default: begin
                            lsu_op = LSU_NOP;
                            illegal_inst = 1;
                        end
                    endcase
                end
            end
            ////////////////////////////////////////////////////////////
            // END: LOAD/STORE Instructions
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: MISC-MEM Instructions
            ////////////////////////////////////////////////////////////
            MISC_MEM: begin
                branch          = 0;
                branch_addr     = 0;
                rs1_en          = 0;
                rs2_en          = 0;
                csr_rd_en       = 0;
                csr_explicit_rd = 0;
                src1            = 0;
                src2            = 0;
                alt_data        = 0;
                alu_op          = ALU_NOP;
                lsu_op          = LSU_NOP;
                case (funct3)
                    FUNCT3_FENCE: begin
                        if (inst[31:28] || rs1_addr || dest_addr) begin // must all be zero
                            illegal_inst = 1;
                        end
                    end
                    FUNCT3_FENCE_I: begin
                        if (inst[31:20] || rs1_addr || dest_addr) begin // must all be zero
                            illegal_inst = 1;
                        end
                    end
                    default: begin
                        illegal_inst = 1;
                    end
                endcase
            end
            ////////////////////////////////////////////////////////////
            // END: MISC-MEM Instructions
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: System Instructions
            ////////////////////////////////////////////////////////////
            SYSTEM: begin
                branch          = 0;
                branch_addr     = 0;
                if (funct3 == 3'b000) begin
                    rs1_en          = 0;
                    rs2_en          = 0;
                    csr_rd_en       = 0;
                    csr_explicit_rd = 0;
                    src1            = 0;
                    src2            = 0;
                    alt_data        = 0;
                    alu_op          = ALU_NOP;
                    lsu_op          = LSU_NOP;
                    if (rs1_addr || dest_addr) begin
                        illegal_inst = 1;
                    end
                    else begin
                        case (funct12)
                            FUNCT12_ECALL:  ecall = 1;
                            FUNCT12_EBREAK: ebreak = 1;
                            FUNCT12_MRET:   mret = 1;
                            FUNCT12_WFI:    ; // NOP
                            default:        illegal_inst = 1;
                        endcase
                    end
                end // if (funct3 == 3'b000)
                else begin
                    // CSR Instructions
                    rs1_en          = (funct3[2]) ? 0 : 1;
                    rs2_en          = 0;
                    csr_rd_en       = 1;
                    csr_explicit_rd = (dest_addr == 0) ? 0 : 1; // explicit read only of destination is not x0
                    src2            = csr_rd_data;
                    alt_data        = csr_rd_data;
                    atomic_csr      = csr_addr_is_atomic & (lsu_op == LSU_CSRRW);
                    illegal_inst    = csr_addr_is_illegal;
                    case (funct3)
                        FUNCT3_CSRRW: begin // read/write
                            src1            = rs1_data;
                            alu_op          = ALU_NOP;
                            lsu_op          = LSU_CSRRW;
                        end
                        FUNCT3_CSRRS: begin // read and set
                            src1            = rs1_data;
                            alu_op          = ALU_OR;
                            lsu_op          = (rs1_addr) ? LSU_CSRRW : LSU_CSRR; // don't write if source is x0
                        end
                        FUNCT3_CSRRC: begin // read and clear
                            src1            = ~rs1_data;
                            alu_op          = ALU_AND;
                            lsu_op          = (rs1_addr) ? LSU_CSRRW : LSU_CSRR; // don't write if source is x0
                        end
                        FUNCT3_CSRRWI: begin // read/write immediate
                            src1            = { {27{1'b0}}, inst[19:15] }; // unsigned, zero-extended
                            alu_op          = ALU_NOP;
                            lsu_op          = LSU_CSRRW;
                        end
                        FUNCT3_CSRRSI: begin // read and set immediate
                            src1            = { {27{1'b0}}, inst[19:15] }; // unsigned, zero-extended
                            alu_op          = ALU_OR;
                            lsu_op          = (inst[19:15]) ? LSU_CSRRW : LSU_CSRR; // don't write if immediate is 0
                        end
                        FUNCT3_CSRRCI: begin // read and clear immediate
                            src1            = ~{ {27{1'b0}}, inst[19:15] }; // unsigned, zero-extended
                            alu_op          = ALU_AND;
                            lsu_op          = (inst[19:15]) ? LSU_CSRRW : LSU_CSRR; // don't write if immediate is 0
                        end
                        default: begin
                            src1    = 0;
                            alu_op  = ALU_NOP;
                            lsu_op  = LSU_NOP;
                            csr_rd_en = 0;
                            csr_explicit_rd = 0;
                            illegal_inst = 1;
                        end
                    endcase
                end
            end
            ////////////////////////////////////////////////////////////
            // END: System Instructions
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: Default (Illegal Instruction)
            ////////////////////////////////////////////////////////////
            default: begin // illegal instruction
                branch = 0;
                branch_addr = 0;
                rs1_en = 0;
                rs2_en = 0;
                csr_rd_en = 0;
                csr_explicit_rd = 0;
                src1 = 0;
                src2 = 0;
                alt_data = 0;
                alu_op = ALU_NOP;
                lsu_op = LSU_NOP;
                illegal_inst = 1;
            end
            ////////////////////////////////////////////////////////////
            // END: Default (Illegal Instruction)
            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////

        endcase
    end

endmodule
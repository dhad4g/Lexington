`timescale 1ns/1ps


module decoder #(
        parameter WIDTH             = 32,               // data width

        localparam OPCODE_WIDTH     = 7,                // RISC-V major opcode width
        localparam REG_ADDR_WIDTH   = 6,                // register file address width
        localparam CSR_ADDR_WIDTH   = 12,               // CSR address width
        localparam ALU_OP_WIDTH     = 4,                // ALU operation select width
        localparam LSU_OP_WIDTH     = 4                 // LSU operation select width
    ) (
        // clock not needed; module is purely combinatorial
        // reset not needed; module is stateless

        input  wire [WIDTH-1:0] inst,                   // instruction bits from fetch
        input  wire [WIDTH-1:0] pc,                     // current program counter
        output wire [WIDTH-1:0] next_pc,                // next PC calculation

        // Register File Ports
        output reg  rs1_en,                             // register source 1 enable
        output wire [REG_ADDR_WIDTH-1:0] rs1_addr,      // register source 1 address
        input  wire [WIDTH-1:0] rs1_data,               // register source 1 data
        output reg  rs2_en,                             // register source 2 enable
        output wire [REG_ADDR_WIDTH-1:0] rs2_addr,      // register source 2 address
        input  wire [WIDTH-1:0] rs2_data,               // register source 2 data

        // CSR Ports
        output reg  csr_rd_en,                          // CSR read enable
        output reg  csr_explicit_rd,                    // CSR explicit read flag
        output wire [CSR_ADDR_WIDTH-1:0] csr_addr,      // CSR read address
        input  wire [WIDTH-1:0] csr_rd_data,            // CSR read data

        // ALU Ports
        output reg  [ALU_OP_WIDTH-1:0] alu_op,          // ALU operation select
        output reg  [WIDTH-1:0] src1,                   // ALU left-side operand
        output reg  [WIDTH-1:0] src2,                   // ALU right-side operand
        input  wire alu_zero                            // ALU zero flag

        // Load/Store Ports
        output reg  [LSU_OP_WIDTH-1:0] lsu_op,          // LSU operation select
        output reg  [WIDTH-1:0] alt_data,               // LSU alternate data
        output wire [REG_ADDR_WIDTH-1:0] dest_addr,     // LSU destination register address
        input  wire dbus_wait,                          // DBus wait signal, suspend until DBus op completes

        // Exception Flags
        output reg  illegal_inst,                       // illegal instruction flag
        output reg  inst_misaligned,                    // instruction misaligned flag, generated by jump/branch instruction
        output reg  ecall,                              // environment call exception flag
        output reg  ebreak,                             // environment breakpoint exception flag
        output reg  mret                                // MRET instruction flag
    );

    // Major OpCode Values
    localparam OP       = 7'b001_0011;
    localparam OP_IMM   = 7'b011_0011;
    localparam LUI      = 7'b011_0111;
    localparam AUIPC    = 7'b001_0111;
    localparam JAL      = 7'b110_1111;
    localparam JALR     = 7'b110_0111;
    localparam BRANCH   = 7'b110_0011;
    localparam LOAD     = 7'b000_0011;
    localparam STORE    = 7'b010_0011;
    localparam MISC_MEM = 7'b000_1111;
    localparam SYSTEM   = 7'b111_0011;

    // Funct7 and Funct3 Field Values
    localparam FUNCT7_ZERO      = 7'b000_0000;
    localparam FUNCT7_BIT30     = 7'b010_0000;
    // arithemetic and logic instructions funct3
    localparam FUNCT3_ADD_SUB   = 3'b000;
    localparam FUNCT3_SHIFT_L   = 3'b001;
    localparam FUNCT3_SLT       = 3'b010;
    localparam FUNCT3_SLTU      = 3'b011;
    localparam FUNCT3_XOR       = 3'b100;
    localparam FUNCT3_SHIFT_R   = 3'b101;
    localparam FUNCT3_OR        = 3'b110;
    localparam FUNCT3_AND       = 3'b111;
    // branch instructions funct3
    localparam FUNCT3_BEQ       = 3'b000;
    localparam FUNCT3_BNE       = 3'b001;
    localparam FUNCT3_BLT       = 3'b100;
    localparam FUNCT3_BGE       = 3'b101;
    localparam FUNCT3_BLTU      = 3'b110;
    localparam FUNCT3_BGEU      = 3'b111;
    // load/store unstruction funct3
    localparam FUNCT3_LB        = 3'b000;
    localparam FUNCT3_LH        = 3'b001;
    localparam FUNCT3_LW        = 3'b010;
    localparam FUNCT3_LBU       = 3'b100;
    localparam FUNCT3_LHU       = 3'b101;
    localparam FUNCT3_SB        = 3'b000;
    localparam FUNCT3_SH        = 3'b001;
    localparam FUNCT3_SW        = 3'b010;
    // fence instruction funct3
    localparam FUNCT3_FENCE     = 3'b000;
    localparam FUNCT3_FENCE_I   = 3'b001;
    // CSR instruction funct3
    localparam FUNCT3_CSRRW     = 3'b001;
    localparam FUNCT3_CSRRS     = 3'b010;
    localparam FUNCT3_CSRRC     = 3'b011;
    localparam FUNCT3_CSRRWI    = 3'b101;
    localparam FUNCT3_CSRRSI    = 3'b110;
    localparam FUNCT3_CSRRCI    = 3'b111;
    // system instructions funct12
    localparam FUNCT12_ECALL    = 12'b0000_0000_0000;
    localparam FUNCT12_EBREAK   = 12'b0000_0000_0001;
    localparam FUNCT12_MRET     = 12'b0011_0000_0010;
    localparam FUNCT12_WFI      = 12'b0001_0000_0101;


    // Internal ALU op select
    localparam ALU_ADD  = 4'b0000;
    localparam ALU_SLL  = 4'b0001;
    localparam ALU_SLTU = 4'b0010;
    localparam ALU_SGEU = 4'b0011;
    localparam ALU_XOR  = 4'b0100;
    localparam ALU_SRL  = 4'b0101;
    localparam ALU_OR   = 4'b0110;
    localparam ALU_AND  = 4'b0111;
    localparam ALU_SUB  = 4'b1000;
    localparam ALU_SLT  = 4'b1010;
    localparam ALU_SGE  = 4'b1011;
    localparam ALU_SRA  = 4'b1101;
    localparam ALU_NOP  = 4'b1111;


    // Internal Load/Store Unit op select
    localparam LSU_LB       = 4'b0000;
    localparam LSU_LH       = 4'b0001;
    localparam LSU_LW       = 4'b0010;
    localparam LSU_LBU      = 4'b0100;
    localparam LSU_LHU      = 4'b0101;
    localparam LSU_SB       = 4'b1000;
    localparam LSU_SH       = 4'b1001;
    localparam LSU_SW       = 4'b1010;
    localparam LSU_CSRR     = 4'b1100;
    localparam LSU_CSRRW    = 4'b1101;
    localparam LSU_REG      = 4'b1110;
    localparam LSU_NOP      = 4'b1111;


    // RISC-V instruction fields
    wire [OPCODE_WIDTH-1:0] opcode;
    wire [REG_ADDR_WIDTH-1:0] dest_addr;
    wire [2:0] funct3;
    wire [6:0] funct7;
    wire [11:0] funct12;
    assign opcode       = inst[6:0];
    assign dest_addr    = inst[11:7];   // output port
    assign funct3       = inst[14:12];
    assign rs1_addr     = inst[19:15];  // output port
    assign rs2_addr     = inst[24:20];  // output port
    assign funct7       = inst[31:25];
    assign funct12      = inst[31:20];
    assign csr_addr     = inst[31:20];  // output port

    // Decode immediate value
    wire [31:0] immediate;
    always_comb begin
        case (opcode)
            OP_IMM:     immediate = { 20{inst[31]}, inst[31:20] }; // sign-extended 12-bit imm[11:0]
            LUI, AUIPC: immediate = { inst[31:12], 12{0}}; // 20-bit upper-immediate imm[31:12], lower bits zero filled
            JAL:        immediate = { 12{inst[31]}, inst[19:12], inst[20], inst[30:21], 0 } // sign-extended 20-bit imm[20:1], lowest bit zeroed
            JAL:        immediate = { 20{inst[31]}, inst[31:20] }; // sign-extended 12-bit imm[11:0]
            BRANCH:     immediate = { 20{inst[31]}, inst[7], inst[30:25], inst[11:8], 0 } // signed-extended 12-bit imm[12:1], lowest bit zeroed
            LOAD:       immediate = { 20{inst[31]}, inst[31:20] }; // sign-extended 12-bit imm[11:0]
            STORE:      immediate = { 20{inst[31]}, inst[31:25], inst[11:7] }; // sign-extended 12-bit imm[11:0]
            MISC-MEM:   immediate = { 20{inst[31]}, inst[31:20] }; // sign-extended 12-bit imm[11:0]
            default:    immediate = { 20{inst[31]}, inst[31:20] }; // most common decoding as default
        endcase
    end

    always_comb begin
        // defaults for exception flags, overwrite per instruction
        inst_misaligned = |(next_pc[1:0]);
        illegal_inst = 0;
        ecall = 0;
        ebreak = 0;
        mret = 0;
        case (opcode)

            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: OP Instructions
            ////////////////////////////////////////////////////////////
            OP: begin
                // Calculate PC
                next_pc = pc + 4;
                // Source read enable
                rs1_en = 1;
                rs2_en = 1;
                csr_rd_en = 0;
                csr_explicit_rd = 0;
                // Source and alt data
                src1 = rs1_data;
                src2 = rs2_data;
                alt_data = 0;
                // LSU OP
                lsu_op = LSU_REG
                // ALU OP
                if (funct7 == FUNCT7_ZERO) begin
                    case (funct3)
                        FUNCT3_ADD_SUB: alu_op = ALU_ADD;
                        FUNCT3_SHIFT_L: alu_op = ALU_SLL;
                        FUNCT3_SLT:     alu_op = ALU_SLT;
                        FUNCT3_SLTU:    alu_op = ALU_SLTU;
                        FUNCT3_XOR:     alu_op = ALU_XOR;
                        FUNCT3_SHIFT_R: alu_op = ALU_SRL;
                        FUNCT3_OR:      alu_op = ALU_OR;
                        FUNCT3_AND:     alu_op = ALU_AND;
                        default: begin
                            alu_op = ALU_NOP;
                            lsu_op = LSU_NOP;
                            illegal_inst = 1;
                        end
                    endcase
                end
                else if (funt7 == FUNCT7_BIT30) begin
                    case (funct3)
                        FUNCT3_ADD_SUB: alu_op = ALU_SUB;
                        FUNCT3_SHIFT_R: alu_op = ALU_SRA;
                        default: begin
                            alu_op = ALU_NOP;
                            lsu_op = LSU_NOP;
                            illegal_inst = 1;
                        end
                    endcase
                end
                else begin
                    alu_op = ALU_NOP;
                    lsu_op = LSU_NOP;
                    illegal_inst = 1;
                end
            end
            ////////////////////////////////////////////////////////////
            // END: OP Instructions
            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: OP-IMM Instructions
            ////////////////////////////////////////////////////////////
            OP_IMM: begin
                next_pc         = pc + 4;
                rs1_en          = 1;
                rs2_en          = 0;
                csr_rd_en       = 0;
                csr_explicit_rd = 0;
                src1            = rs1_data;
                src2            = immediate;
                alt_data        = 0;
                lsu_op          = LSU_REG;
                // ALU OP
                if (funct7 == FUNCT7_ZERO) begin
                    case (funct3)
                        FUNCT3_ADD_SUB: alu_op = ALU_ADD;
                        FUNCT3_SHIFT_L: alu_op = ALU_SLL;
                        FUNCT3_SLT:     alu_op = ALU_SLT;
                        FUNCT3_SLTU:    alu_op = ALU_SLTU;
                        FUNCT3_XOR:     alu_op = ALU_XOR;
                        FUNCT3_SHIFT_R: alu_op = ALU_SRL;
                        FUNCT3_OR:      alu_op = ALU_OR;
                        FUNCT3_AND:     alu_op = ALU_AND;
                        default:
                            begin
                                alu_op = ALU_NOP;
                                lsu_op = LSU_NOP;
                                illegal_inst = 1;
                            end
                    endcase
                end
                else if (funt7 == FUNCT7_BIT30) begin
                    case (funct3)
                        FUNCT3_SHIFT_R: alu_op = ALU_SRA;
                        default:
                            begin
                                alu_op = ALU_NOP;
                                lsu_op = LSU_NOP;
                                illegal_inst = 1;
                            end
                    endcase
                end
                else begin
                    alu_op = ALU_NOP;
                    lsu_op = LSU_NOP;
                    illegal_inst = 1;
                end
            end
            ////////////////////////////////////////////////////////////
            // END: OP-IMM Instructions
            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: LUI/AUIPC Instructions
            ////////////////////////////////////////////////////////////
            LUI, AUIPC: begin
                next_pc         = pc + 4;
                rs1_en          = 0;
                rs2_en          = 0;
                csr_rd_en       = 0;
                csr_explicit_rd = 0;
                src1            = (opcode == AUIPC) ? pc : 0;
                src2            = immediate;
                alt_data        = 0;
                alu_op          = ALU_ADD;
                lsu_op          = LSU_REG;
            end
            ////////////////////////////////////////////////////////////
            // END: LUI/AUIPC Instructions
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: JAL/JALR Instruction
            ////////////////////////////////////////////////////////////
            JAL, JALR: begin
                rs1_en          = (opcode == JALR) ? 1 : 0;
                rs2_en          = 0;
                csr_rd_en       = 0;
                csr_explicit_rd = 0;
                src1            = pc;
                src2            = 4;
                alt_data        = 0;
                alu_op          = ALU_ADD;
                lsu_op          = LSU_REG;
                // calculate jump address
                if (opcode == JAL) begin
                    next_pc     = pc + immediate;
                end
                else begin // JALR
                    // sign-extended immediate, lowet bit zeroed after calculation
                    next_pc[31:1] = (rs1_data + immediate)[31:1];
                    next_pc[0]    = 0;
                end
                if (inst_misaligned) begin
                    lsu_op = LSU_NOP;
                end
            end
            ////////////////////////////////////////////////////////////
            // END: JAL/JALR Instruction
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: BRANCH Instructions
            ////////////////////////////////////////////////////////////
            BRANCH: begin
                rs1_en          = 1;
                rs2_en          = 1;
                csr_rd_en       = 0;
                csr_explicit_rd = 0;
                src1            = rs1_data;
                src2            = rs2_data;
                alt_data        = 0;
                lsu_op          = LSU_NOP;
                // Next PC
                // sign-extended immediate, lowest bit zero
                if (funct3 == FUNCT3_BEQ) begin
                    next_pc     = (alu_zero)  ? (pc + immediate) : (pc + 4);
                end
                else begin
                    next_pc     = (!alu_zero) ? (pc + immediate) : (pc + 4);
                end
                // ALU OP
                case (funct3)
                    FUNCT3_BEQ:     alu_op = ALU_XOR;  // branch if equal
                    FUNCT3_BNE:     alu_op = ALU_XOR;  // branch if not equal
                    FUNCT3_BLT:     alu_op = ALU_SLT;  // branch if less than
                    FUNCT3_BGE:     alu_op = ALU_SGE;  // branch if greater than or equal
                    FUNCT3_BLTU:    alu_op = ALU_SLTU: // branch if less than unsigned
                    FUNCT3_BGEU:    alu_op = ALU_SGEU: // branch if greater than or equal unsigned
                    default: begin
                        alu_op  = ALU_NOP;
                        illegal_inst = 1;
                    end
                endcase
            end
            ////////////////////////////////////////////////////////////
            // END: BRANCH Instructions
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: LOAD/STORE Instuctions
            ////////////////////////////////////////////////////////////
            LOAD, STORE: begin
                next_pc         = pc + 4;
                rs1_en          = 1;
                rs2_en          = (opcode == STORE) ? 1 : 0;
                csr_rd_en       = 0;
                csr_explicit_rd = 0;
                src1            = rs1_data;
                src2            = immediate;
                alt_data        = (opcode == STORE) ? rs2_data : 0;
                alu_op          = ALU_ADD;
                if (opcode == LOAD) begin
                    case (funct3)
                        FUNCT3_LB:  lsu_op = LSU_LB;
                        FUNCT3_LH:  lsu_op = LSU_LH;
                        FUNCT3_LW:  lsu_op = LSU_LW;
                        FUNCT3_LBU: lsu_op = LSU_LBU;
                        FUNCT3_LHU: lsu_op = LSU_LHU;
                        default: begin
                            lsu_op = LSU_NOP;
                            illegal_inst = 1;
                        end
                    endcase
                end
                else begin // STORE
                    case (funct3)
                        FUNCT3_SB:  lsu_op = LSU_SB;
                        FUNCT3_SH:  lsu_op = LSU_SH;
                        FUNCT3_SW:  lsu_op = LSU_SW;
                        default: begin
                            lsu_op = LSU_NOP;
                            illegal_inst = 1;
                        end
                    endcase
                end
            end
            ////////////////////////////////////////////////////////////
            // END: LOAD/STORE Instuctions
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: MISC-MEM Instructions
            ////////////////////////////////////////////////////////////
            MISC_MEM: begin
                next_pc         = pc + 4;
                rs1_en          = 0;
                rs2_en          = 0;
                csr_rd_en       = 0;
                csr_explicit_rd = 0;
                src1            = 0;
                src2            = 0;
                alt_data        = 0;
                alu_op          = ALU_NOP;
                lsu_op          = LSU_NOP;
                case (funct3)
                    FUNCT3_FENCE: begin
                        if (inst[31:28] || rs1_addr || dest_addr) begin // must all be zero
                            illegal_inst = 1;
                        end
                    end
                    FUNCT3_FENCE_I: begin
                        if (inst[31:20] || rs1_addr || dest_addr) begin // must all be zero
                            illegal_inst = 1;
                        end
                    end
                    default: begin
                        illegal_inst = 1;
                    end
                endcase
            end
            ////////////////////////////////////////////////////////////
            // END: MISC-MEM Instructions
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: System Instructions
            ////////////////////////////////////////////////////////////
            SYSTEM: begin
                next_pc         = pc + 4;
                if (funct3 == 3'b000) begin
                    rs1_en          = 0;
                    rs2_en          = 0;
                    csr_rd_en       = 0;
                    csr_explicit_rd = 0;
                    src1            = 0;
                    src2            = 0;
                    alt_data        = 0;
                    alu_op          = ALU_NOP;
                    lsu_op          = LSU_NOP;
                    if (rs1_addr || dest_addr) begin
                        illegal_inst = 1;
                    end
                    else begin
                        case (funct12)
                            FUNCT12_ECALL:  ecall = 1;
                            FUNCT12_EBREAK: ebreak = 1;
                            FUNCT12_MRET:   mret = 1;
                            FUNCT12_WFI:    ; // NOP
                            default:        illegal_inst = 1;
                        endcase
                    end
                end
                else begin
                    // CSR Instructions
                    rs1_en          = (funct3[2]) ? 0 : 1;
                    rs2_en          = 0;
                    csr_rd_en       = 1;
                    csr_explicit_rd = (dest_addr == 0) ? 0 : 1; // explicit read only of destination is not x0
                    src2            = csr_rd_data;
                    alt_data        = csr_rd_data;
                    case (funct3)
                        FUNCT3_CSRRW: begin // read/write
                            src1            = rs1_data;
                            alu_op          = ALU_NOP;
                            lsu_op          = LSU_CSRRW;
                        end
                        FUNCT3_CSRRS: begin // read and set
                            src1            = rs1_data;
                            alu_op          = ALU_OR;
                            lsu_op          = (rs1_addr) ? LSU_CSRRW : LSU_CSRR; // don't write if source is x0
                        end
                        FUNCT3_CSRRC: begin // read and clear
                            src1            = ~rs1_data;
                            alu_op          = ALU_AND;
                            lsu_op          = (rs1_addr) ? LSU_CSRRW : LSU_CSRR; // don't write if source is x0
                        end
                        FUNCT3_CSRRWI: begin // read/write immediate
                            src1            = { 27{0}, inst[19:15] }; // unsigned, zero-extended
                            alu_op          = ALU_NOP;
                            lsu_op          = LSU_CSRRW;
                        end
                        FUNCT3_CSRRSI: begin // read and set immediate
                            src1            = { 27{0}, inst[19:15] }; // unsigned, zero-extended
                            alu_op          = ALU_OR;
                            lsu_op          = (inst[19:15]) ? LSU_CSRRW : LSU_CSRR; // don't write if immediate is 0
                        end
                        FUNCT3_CSRRCI: begin // read and clear immediate
                            src1            = ~{ 27{0}, inst[19:15] }; // unsigned, zero-extended
                            alu_op          = ALU_AND;
                            lsu_op          = (inst[19:15]) ? LSU_CSRRW : LSU_CSRR; // don't write if immediate is 0
                        end
                        default: begin
                            src1    = 0;
                            alu_op  = ALU_NOP;
                            lsu_OP  = LSU_NOP;
                            csr_rd_en = 0;
                            csr_explicit_rd = 0;
                            illegal_inst = 1;
                        end
                    endcase
                end
            end
            ////////////////////////////////////////////////////////////
            // END: System Instructions
            ////////////////////////////////////////////////////////////


            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////
            // BEGIN: Default (Illegal Instruction)
            ////////////////////////////////////////////////////////////
            default: begin // illegal instruction
                next_pc = pc + 4;
                rs1_en = 0;
                rs2_en = 0;
                csr_rd_en = 0;
                csr_explicit_rd = 0;
                src1 = 0;
                src2 = 0;
                alt_data = 0;
                alu_op = ALU_NOP;
                lsu_op = LSU_NOP;
                illegal_inst = 1;
            end
            ////////////////////////////////////////////////////////////
            // END: Default (Illegal Instruction)
            ////////////////////////////////////////////////////////////
            ////////////////////////////////////////////////////////////

        endcase
    end

endmodule
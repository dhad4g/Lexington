`ifndef __AXI4_LITE_SV
`define __AXI4_LITE_SV


interface axi4_lite #(
        parameter WIDTH         = 32,       // data bus width
        parameter ADDR_WIDTH    = 32        // address bus width
    );

        typedef struct packed {
            logic privileged;
            logic non_secure;
            logic inst_data_n;
        } prot_t;

        typedef enum logic [1:0] {
            OKAY    = 2'b00,
            EXOKAY  = 2'b01,    // exclusive access okay, invalid for AXI4-Lite
            SLVERR  = 2'b10,    // subordinate error
            DECERR  = 2'b11     // decode error, generated by interconnect
        } resp_t;

        // Global signals
        logic aclk;
        logic areset_n;
        // Write address channel
        logic awvalid;
        logic awready;
        logic [ADDR_WIDTH-1:0] awaddr;
        prot_t awprot;
        // Write data channel
        logic wvalid;
        logic wready;
        logic [WIDTH-1:0] wdata;
        logic [(WIDTH/8)-1:0] wstrb;
        // Write response channel
        logic bvalid;
        logic bready;
        resp_t bresp;
        // Read address channel
        logic arvalid;
        logic arready;
        logic [ADDR_WIDTH-1:0] araddr;
        prot_t arprot;
        // Read data channel
        logic rvalid;
        logic rready;
        logic [WIDTH-1:0] rdata;
        resp_t rresp;


        modport manager (
            output aclk, output areset_n, // global signals
            output awvalid, input  awready, output awaddr, output awprot, // write address channel
            output wvalid, input  wready, output wdata, output wstrb, // write data channel
            input  bvalid, output bready, input  bresp, // write response channel
            output arvalid, input  arready, output araddr, output arprot, // read address channel
            input  rvalid, output rready, input  rdata, input rresp // read data channel
        );

        modport subordinate (
            input aclk, input areset_n, // global signals
            input awvalid, output  awready, input awaddr, input awprot, // write address channel
            input wvalid, output  wready, input wdata, input wstrb, // write data channel
            output  bvalid, input bready, output  bresp, // write response channel
            input arvalid, output  arready, input araddr, input arprot, // read address channel
            output  rvalid, input rready, output  rdata, output rresp // read data channel
        );

endinterface

`endif //__AXI4_LITE_SV
`timescale 1ns/1ps

`include "rv32.sv"
`include "lexington.sv"
import lexington::*;


module dbus #(
        parameter ROM_ADDR_WIDTH    = DEFAULT_ROM_ADDR_WIDTH,       // ROM address width (word-addressable, default 4kB)
        parameter RAM_ADDR_WIDTH    = DEFAULT_RAM_ADDR_WIDTH,       // RAM address width (word-addressable, default 4kB)
        localparam MTIME_ADDR_WIDTH = 2,
        parameter AXI_ADDR_WIDTH    = DEFAULT_AXI_ADDR_WIDTH,       // AXI bus address space width (byte-addressable)
        parameter ROM_BASE_ADDR     = DEFAULT_ROM_BASE_ADDR,        // ROM base address (must be aligned to ROM size)
        parameter RAM_BASE_ADDR     = DEFAULT_RAM_BASE_ADDR,        // RAM base address (must be aligned to RAM size)
        parameter MTIME_BASE_ADDR   = DEFAULT_MTIME_BASE_ADDR,      // machine timer base address (see [CSR](./CSR.md))
        parameter AXI_BASE_ADDR     = DEFAULT_AXI_BASE_ADDR        // AXI bus address space base (must be aligned to AXI address space)
    ) (
        // clock not needed; module is asynchronous
        // reset not needed; module is read-only

        input  logic rd_en,                                         // read enable from LSU
        input  logic wr_en,                                         // write enable from LSU
        input  rv32::word addr,                                     // read/write address from LSU
        input  rv32::word wr_data_i,                                // write data from LSU
        input  logic [(rv32::XLEN/8)-1:0] wr_strobe_i,              // write strobe (input)
        input  rv32::word rom_rd_data,                              // read data from ROM
        input  rv32::word ram_rd_data,                              // read data from RAM
        input  rv32::word mtime_rd_data,                            // read data from mtime module
        input  rv32::word axi_rd_data,                              // read data from AXI interface
        input  logic axi_access_fault,                              // flag indicating AXI transaction access fault
        input  logic axi_busy,                                      // flag indicating AXI transaction requires additonal cycles

        output rv32::word rd_data,                                  // read data to LSU
        output logic rom_rd_en,                                     // read enable to ROM
        output logic [ROM_ADDR_WIDTH-1:0] rom_addr,                 // *word-addressable* address to ROM
        output logic ram_rd_en,                                     // read enable to RAM
        output logic ram_wr_en,                                     // write enable to RAM
        output logic [RAM_ADDR_WIDTH-1:0] ram_addr,                 // *word-addressable* address to RAM
        output logic mtime_rd_en,                                   // read enable to mtime module
        output logic mtime_wr_en,                                   // write enable to mtime module
        output logic [MTIME_ADDR_WIDTH-1:0] mtime_addr,             // *word-addressable* address to mtime module
        output logic axi_rd_en,                                     // read enable to AXI interface
        output logic axi_wr_en,                                     // write enable to AXI interface
        output logic [AXI_ADDR_WIDTH-1:0] axi_addr,                 // *byte-addressable* address to AXI interface
        output rv32::word wr_data_o,                                // shared write data to ROM/RAM/mtime/AXI
        output logic [(rv32::XLEN/8)-1:0] wr_strobe_o,              // write strobe (output)
        output logic data_misaligned,                               // asserted if memory address is not 4-byte aligned
        output logic data_access_fault,                             // access fault flag to Trap Unit
        output logic load_store_n,                                  // indicates if exception was generated by load or store(0=store,1=load)
        output logic dbus_wait,                                     // asserted if dbus transaction requires additional cycles
        output logic dbus_err                                       // logical or of data_misaligned and data_access_fault
    );

    // Address space mask function
    function automatic rv32::word mask_upper_bits(rv32::word addr, integer bit_width);
        rv32::word mask;
        mask = (~(0)) << bit_width;
        return mask & addr;
    endfunction


    // Word-addressable address
    localparam WORD_ADDR_WIDTH = rv32::XLEN - rv32::ADDR_BITS_IN_WORD;
    logic [WORD_ADDR_WIDTH-1:0] word_addr;
    assign word_addr = addr >> rv32::ADDR_BITS_IN_WORD;

    // Select address bits
    assign rom_addr     = word_addr[ROM_ADDR_WIDTH-1:0];        // word-addressable
    assign ram_addr     = word_addr[RAM_ADDR_WIDTH-1:0];        // word-addressable
    assign mtime_addr   = word_addr[MTIME_ADDR_WIDTH-1:0];      // word-addressable
    assign axi_addr     = addr[AXI_ADDR_WIDTH-1:0];             // byte-addressable

    // Detect address space
    logic is_rom_addr, is_ram_addr, is_mtime_addr, is_axi_addr;
    assign is_rom_addr      = (ROM_BASE_ADDR == mask_upper_bits(addr, ROM_ADDR_WIDTH + rv32::ADDR_BITS_IN_WORD));       // word-addressable
    assign is_ram_addr      = (RAM_BASE_ADDR == mask_upper_bits(addr, RAM_ADDR_WIDTH + rv32::ADDR_BITS_IN_WORD));       // word-addressable
    assign is_mtime_addr    = (MTIME_BASE_ADDR == mask_upper_bits(addr, MTIME_ADDR_WIDTH + rv32::ADDR_BITS_IN_WORD));   // word-addressable
    assign is_axi_addr      = (AXI_BASE_ADDR == mask_upper_bits(addr, AXI_ADDR_WIDTH));                                 // byte-addressable


    // Set data_misaligned, load_store_n, and dbus_wait
    assign data_misaligned  = (rd_en | wr_en) & (|(addr[rv32::ADDR_BITS_IN_WORD-1:0]));
    assign load_store_n     = rd_en;
    assign dbus_wait        = ((rd_en | wr_en) && is_axi_addr) ? axi_busy : 0;
    assign dbus_err         = data_misaligned | data_access_fault;

    // Pass through wr_data and wr_strobe
    assign wr_data_o = wr_data_i;
    assign wr_strobe_o = wr_strobe_i;

    // Read/Write enable and read data routing
    always_comb begin
        // default data_access_fault to 0
        data_access_fault = 0;
        // default all rd/wr enable to 0
        rom_rd_en = 0;
        ram_rd_en = 0;
        ram_wr_en = 0;
        mtime_rd_en = 0;
        mtime_wr_en = 0;
        axi_rd_en = 0;
        axi_wr_en = 0;
        rd_data   = 0;
        if (!data_misaligned) begin
            if (is_rom_addr) begin
                if (wr_en) begin // write permission prohibited
                    data_access_fault = 1;
                    rd_data = 0;
                end
                else begin
                    rom_rd_en = rd_en;
                    rd_data   = rom_rd_data;
                end
            end
            else if (is_ram_addr) begin
                ram_rd_en = rd_en;
                ram_wr_en = wr_en;
                rd_data = ram_rd_data;
            end
            else if (is_mtime_addr) begin
                mtime_rd_en = rd_en;
                mtime_wr_en = wr_en;
                rd_data = mtime_rd_data;
            end
            else if (is_axi_addr) begin
                data_access_fault = axi_access_fault;
                axi_rd_en = rd_en;
                axi_wr_en = wr_en;
                rd_data = axi_rd_data;
            end
            else begin
                data_access_fault = rd_en | wr_en;
                rd_data = 0;
            end
        end // if (!data_misaligned)
    end


endmodule

`timescale  1ns/1ps

`include rv32.sv
`include saratoga.sv


module control (
        input  logic clk,
        input  logic rst_n,
    );

endmodule
